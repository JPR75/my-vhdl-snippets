-------------------------------------------------------------------------------
-- Title   : Constant
-- Project : Digilent X3S1600E eval board test
-------------------------------------------------------------------------------
-- Description : Constant declaration
-------------------------------------------------------------------------------
-- File     : const.vhdl
-- Revision : 1.0.0
-- Created  : April 24, 2011
-- Updated  : April 24, 2011
-------------------------------------------------------------------------------
-- Author       : JPR75
-- Web          : -
-- Email        : -
-------------------------------------------------------------------------------
-- Licence : GNU GPL
--           -
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
package const is

  constant c_CLK_50MHz : real := 50000000.0; -- 50MHz on board CLK

end const;

-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
package body const is


end package body const;

